module top_module(inputa, input b, output c);
assign y= a&b;
endmodule

